module FSM(
  input In1,
  input RST,
  input CLK, 
  output reg Out1
);
reg [1:0] state;
	
	// Declare states
	parameter S0 = 0, S1 = 1, S2 = 2, S3 = 3;
	
	// Output depends only on the state
	always @ (state) begin
		case (state)
			S0:
				Out1 = 2'b01;
			S1:
				Out1 = 2'b10;
			S2:
				Out1 = 2'b11;
			S3:
				Out1 = 2'b00;
			default:
				Out1 = 2'b00;
		endcase
	end
	
	// Determine the next state
	always @ (posedge CLK or posedge RST) begin
		if (RST)
			state <= S0;
		else
			case (state)
				S0:
					state <= S1;
				S1:
					if (In1)
						state <= S2;
					else
						state <= S1;
				S2:
					if (In1)
						state <= S3;
					else
						state <= S1;
				S3:
					if (In1)
						state <= S2;
					else
						state <= S3;
			endcase
	end

endmodule 